/* synthesis translate_off*/
`define SBP_SIMULATION
/* synthesis translate_on*/
`ifndef SBP_SIMULATION
`define SBP_SYNTHESIS
`endif

//
// Verific Verilog Description of module FIFO_buffer
//
module FIFO_buffer () /* synthesis sbp_module=true */ ;
    
    
    fifo_16bit fifo_16bit_inst ();
    
endmodule

