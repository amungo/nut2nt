--VHDL instantiation template

component FIFO_buffer is
    
end component FIFO_buffer; -- sbp_module=true 
_inst: FIFO_buffer port map ();
