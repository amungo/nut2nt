/* synthesis translate_off*/
`define SBP_SIMULATION
/* synthesis translate_on*/
`ifndef SBP_SIMULATION
`define SBP_SYNTHESIS
`endif

//
// Verific Verilog Description of module FIFO_buffer
//
module FIFO_buffer () /* synthesis sbp_module=true */ ;
    
    
    fifo_8bit_buffer fifo_8bit_buffer_inst ();
    fifo_8bit_sl fifo_8bit_sl_inst ();
    
endmodule

